// Nios2Computer_tb.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module Nios2Computer_tb (
	);

	wire        nios2computer_inst_clk_bfm_clk_clk;               // Nios2Computer_inst_clk_bfm:clk -> [Nios2Computer_inst:clk_clk, Nios2Computer_inst_reset_bfm:clk]
	wire  [7:0] nios2computer_inst_led_pio_ext_connection_export; // Nios2Computer_inst:led_pio_ext_connection_export -> Nios2Computer_inst_led_pio_ext_connection_bfm:sig_export
	wire        nios2computer_inst_reset_bfm_reset_reset;         // Nios2Computer_inst_reset_bfm:reset -> Nios2Computer_inst:reset_reset_n

	Nios2Computer nios2computer_inst (
		.clk_clk                       (nios2computer_inst_clk_bfm_clk_clk),               //                    clk.clk
		.led_pio_ext_connection_export (nios2computer_inst_led_pio_ext_connection_export), // led_pio_ext_connection.export
		.reset_reset_n                 (nios2computer_inst_reset_bfm_reset_reset)          //                  reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios2computer_inst_clk_bfm (
		.clk (nios2computer_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm nios2computer_inst_led_pio_ext_connection_bfm (
		.sig_export (nios2computer_inst_led_pio_ext_connection_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) nios2computer_inst_reset_bfm (
		.reset (nios2computer_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (nios2computer_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
